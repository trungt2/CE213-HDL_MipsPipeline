library verilog;
use verilog.vl_types.all;
entity tb_cpu is
end tb_cpu;
